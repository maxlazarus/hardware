CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 130 30 100 9
0 68 1366 418
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 68 1366 418
1217921043 0
0
6 Title:
5 Name:
0
0
0
14
10 P-EMOS 3T~
219 405 284 0 3 7
0 3 12 10
0
0 0 848 692
7 IRF9510
17 0 66 8
2 Q1
35 -10 49 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-220
7

0 2 1 3 2 1 3 0
109 0 0 256 1 0 0 0
1 Q
8953 0 0
0
0
10 P-EMOS 3T~
219 311 286 0 3 7
0 3 8 11
0
0 0 848 692
7 IRF9510
17 0 66 8
2 Q4
35 -10 49 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-220
7

0 2 1 3 2 1 3 0
109 0 0 256 1 0 0 0
1 Q
4441 0 0
0
0
10 N-EMOS 3T~
219 533 320 0 3 7
0 6 3 7
0
0 0 848 0
9 IRFI1010G
17 0 80 8
2 Q3
42 -10 56 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-220
7

0 2 3 1 2 3 1 0
77 0 0 256 1 0 0 0
1 Q
3618 0 0
0
0
10 N-EMOS 3T~
219 676 320 0 3 7
0 5 4 7
0
0 0 848 0
9 IRFI1010G
17 0 80 8
2 Q5
42 -10 56 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-220
7

0 2 3 1 2 3 1 0
77 0 0 256 1 0 0 0
1 Q
6153 0 0
0
0
2 +V
167 598 228 0 1 3
0 4
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
2 +V
167 411 241 0 1 3
0 10
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
2 +V
167 206 201 0 1 3
0 9
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 344 391 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
2 +V
167 318 240 0 1 3
0 11
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3549 0 0
0
0
2 +V
167 352 200 0 1 3
0 12
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7931 0 0
0
0
9 Resistor~
219 682 273 0 4 5
0 5 4 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 538 272 0 3 5
0 4 6 1
0
0 0 880 270
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 207 255 0 4 5
0 8 9 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 344 343 0 3 5
0 2 3 -1
0
0 0 880 90
4 100k
2 0 30 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
16
0 2 3 0 0 8320 0 0 3 16 0 3
379 303
379 329
515 329
2 0 4 0 0 12416 0 4 0 0 3 4
658 329
658 330
641 330
641 237
1 2 4 0 0 128 0 5 11 0 0 3
598 237
682 237
682 255
1 1 4 0 0 128 0 12 5 0 0 3
538 254
538 237
598 237
1 1 5 0 0 12416 0 4 11 0 0 4
682 302
682 303
682 303
682 291
2 1 6 0 0 8320 0 12 3 0 0 3
538 290
539 290
539 302
0 3 7 0 0 4096 0 0 4 8 0 4
537 372
683 372
683 338
682 338
0 3 7 0 0 4224 0 0 3 0 0 3
344 372
539 372
539 338
1 2 8 0 0 4224 0 13 2 0 0 5
207 273
207 372
262 372
262 277
293 277
1 2 9 0 0 8320 0 7 13 0 0 3
206 210
207 210
207 237
1 3 10 0 0 8320 0 6 1 0 0 4
411 250
412 250
412 266
411 266
1 3 11 0 0 8320 0 9 2 0 0 3
318 249
317 249
317 268
2 1 12 0 0 12416 0 1 10 0 0 6
387 275
387 276
366 276
366 235
352 235
352 209
1 1 2 0 0 4224 0 14 8 0 0 2
344 361
344 385
2 0 3 0 0 0 0 14 0 0 16 2
344 325
344 303
1 1 3 0 0 128 0 2 1 0 0 4
317 304
317 303
411 303
411 302
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2360684 1210432 100 100 0 0
0 0 0 0
0 96 161 166
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2425856 8550464 100 100 0 0
77 66 1337 276
0 418 1366 768
1337 66
77 66
1337 68
1337 276
0 0
5e-006 0 5 5 5e-006 5e-006
12401 0
4 1e-006 2
1
539 296
0 6 0 0 2	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
