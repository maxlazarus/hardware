CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
34 95 1332 751
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
34 95 1332 751
1217921042 0
0
6 Title:
5 Name:
0
0
0
6
7 Ground~
168 580 428 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
9 V Source~
197 798 237 0 2 5
0 3 2
0
0 0 17264 0
2 5V
16 0 30 8
3 Vs2
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
4441 0 0
0
0
9 V Source~
197 376 227 0 2 5
0 5 2
0
0 0 17264 0
2 3V
16 0 30 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3618 0 0
0
0
10 N-EMOS 3T~
219 546 284 0 3 7
0 3 5 4
0
0 0 848 270
4 NMOS
-16 30 12 38
2 Q1
-9 20 5 28
0
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
77 0 0 0 0 0 0 0
1 Q
6153 0 0
0
0
9 Resistor~
219 661 228 0 2 5
0 3 3
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 456 221 0 2 5
0 4 5
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
8
0 0 3 0 0 8192 0 0 0 7 6 3
660 292
736 292
736 178
1 3 4 0 0 8320 0 6 4 0 0 3
456 239
456 292
526 292
0 2 5 0 0 8320 0 0 4 8 0 3
456 179
535 179
535 268
1 0 2 0 0 4096 0 1 0 0 5 2
580 422
580 392
2 2 2 0 0 8320 0 2 3 0 0 4
798 258
798 392
376 392
376 248
2 1 3 0 0 8320 0 5 2 0 0 4
661 210
661 178
798 178
798 216
1 1 3 0 0 128 0 4 5 0 0 3
562 292
661 292
661 246
2 1 5 0 0 128 0 6 3 0 0 4
456 203
456 177
376 177
376 206
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
