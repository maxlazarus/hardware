CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
350 140 30 200 9
5 73 649 763
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
5 73 649 763
1285029907 256
0
6 Title:
5 Name:
0
0
0
15
10 Capacitor~
219 526 378 0 2 5
0 2 5
0
0 0 848 90
3 1uF
11 0 32 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
7 Ground~
168 479 408 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
11 Signal Gen~
195 429 368 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1259902592 0 1041865114
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 704006255
20
1 1e+007 0 0.15 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -150m/150mV
-39 -30 38 -22
2 V3
-7 -40 7 -32
0
0
42 %D %1 %2 DC 0 SIN(0 150m 10Meg 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
10 Capacitor~
219 628 272 0 2 5
0 2 3
0
0 0 848 90
4 10nF
8 0 36 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
2 +V
167 552 260 0 1 3
0 7
0
0 0 54256 0
6 2.048V
-21 -22 21 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
7 Op Amp~
219 510 236 0 3 7
0 8 10 4
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 0 0 0 0
1 U
7734 0 0
0
0
7 Ground~
168 416 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 444 302 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
11 Signal Gen~
195 382 246 0 19 64
0 9 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1259902592 0 1041865114
20
1 1e+007 0 0.15 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -150m/150mV
-39 -30 38 -22
2 V2
-7 -40 7 -32
0
0
42 %D %1 %2 DC 0 SIN(0 150m 10Meg 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3549 0 0
0
0
9 Resistor~
219 600 234 0 2 5
0 4 3
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 494 348 0 2 5
0 6 5
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 506 270 0 3 5
0 7 8 1
0
0 0 880 180
3 10k
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 456 242 0 2 5
0 9 8
0
0 0 880 0
2 1k
-11 16 3 24
2 R4
-9 8 5 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 460 230 0 3 5
0 2 10 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 528 162 0 2 5
0 10 4
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
16
2 2 3 0 0 8320 0 10 4 0 0 3
618 234
628 234
628 263
1 0 4 0 0 4096 0 10 0 0 15 2
582 234
576 234
2 2 5 0 0 4224 0 1 11 0 0 3
526 369
526 348
512 348
1 1 2 0 0 4096 0 2 1 0 0 3
479 402
526 402
526 387
2 1 2 0 0 0 0 3 2 0 0 3
460 373
460 402
479 402
1 1 6 0 0 8320 0 3 11 0 0 3
460 363
460 348
476 348
1 1 2 0 0 16528 0 4 8 0 0 5
628 281
628 295
578 295
578 296
444 296
1 1 7 0 0 4224 0 12 5 0 0 3
524 270
552 270
552 269
0 2 8 0 0 4224 0 0 12 10 0 3
484 242
484 270
488 270
2 1 8 0 0 128 0 13 6 0 0 2
474 242
492 242
1 1 9 0 0 8320 0 13 9 0 0 3
438 242
438 241
413 241
0 1 10 0 0 4224 0 0 15 13 0 3
484 230
484 162
510 162
2 2 10 0 0 128 0 6 14 0 0 2
492 230
478 230
1 1 2 0 0 128 0 14 7 0 0 4
442 230
442 185
416 185
416 184
2 3 4 0 0 8320 0 15 6 0 0 5
546 162
576 162
576 235
528 235
528 236
2 1 2 0 0 128 0 9 8 0 0 3
413 251
413 296
444 296
0
0
2073 0 1
0
0
0
0.1 0.2 0
0
0 0 0
100 2 1 1e+008
0 5e-007 2e-009 2e-009
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
7210002 1210432 100 100 0 0
0 0 0 0
5 73 166 143
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 1
0
4066420 8550976 100 100 0 0
77 66 677 276
637 408 1355 753
677 66
77 66
677 70
677 276
0 0
5e-007 0 3.53143 0 5e-007 5e-007
12409 3
4 1e-007 5
1
577 234
0 4 0 0 1	0 2 0 0
3540154 4421696 100 100 0 0
77 66 669 276
651 69 1346 414
668 66
77 66
669 66
669 276
0 0
9.69363e+007 1 20.299 19.699 9.96247e+007 9.96247e+007
12387 0
4 3e+007 5e+007
1
579 234
0 4 0 0 1	0 2 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
